* Simple hysteresis placeholder
V1 in 0 DC 5
R1 in out 2
C1 out 0 0.02
.tran 0.01 1
.control
run
quit
.endc
.end